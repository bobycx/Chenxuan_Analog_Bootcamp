** sch_path: /mnt/c/Users/ycx/dev/Analog/Chenxuan_Analog_Bootcamp/analog/schematics/bootcamp_opamp.sch
**.subckt bootcamp_opamp
XM1 net2 net1 GND GND sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29' pd='2*int((nf+1)/2) * (W/nf + 0.29)'
+ ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W' sa=0 sb=0 sd=0 mult=1 m=1
V1 net1 GND 0
V2 net2 GND 0.9
**** begin user architecture code



.lib ~/.volare/volare/sky130/versions/fa87f8f4bbcc7255b6f0c0fb506960f531ae2392/sky130B/libs.tech/ngspice/sky130.lib.spice tt

.control
	dc V1 0 3 0.01
	plot -i(V2)

.endc

.save all



**** end user architecture code
**.ends
.GLOBAL GND
.end
